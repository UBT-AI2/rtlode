// addsubfp_single.v

// Generated using ACDS version 17.1.1 273

`timescale 1 ps / 1 ps
module addsubfp_single (
		input  wire [31:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire [31:0] b,      //      b.b
		input  wire        clk,    //    clk.clk
		input  wire [0:0]  opSel,  //  opSel.opSel
		output wire [31:0] q       //      q.q
	);

	addsubfp_single_altera_fp_functions_171_cvdbjfi fp_functions_0 (
		.clk    (clk),    //   input,   width = 1,    clk.clk
		.areset (areset), //   input,   width = 1, areset.reset
		.a      (a),      //   input,  width = 32,      a.a
		.b      (b),      //   input,  width = 32,      b.b
		.q      (q),      //  output,  width = 32,      q.q
		.opSel  (opSel)   //   input,   width = 1,  opSel.opSel
	);

endmodule
