// multfp_double.v

// Generated using ACDS version 17.1.1 273

`timescale 1 ps / 1 ps
module multfp_double (
		input  wire [63:0] a,      //      a.a
		input  wire        areset, // areset.reset
		input  wire [63:0] b,      //      b.b
		input  wire        clk,    //    clk.clk
		output wire [63:0] q       //      q.q
	);

	multfp_double_altera_fp_functions_171_s7r74ky fp_functions_0 (
		.clk    (clk),    //   input,   width = 1,    clk.clk
		.areset (areset), //   input,   width = 1, areset.reset
		.a      (a),      //   input,  width = 64,      a.a
		.b      (b),      //   input,  width = 64,      b.b
		.q      (q)       //  output,  width = 64,      q.q
	);

endmodule
